-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Sat Nov 04 13:00:33 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY AffichagePorte IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        X : IN STD_LOGIC := '0';
        HEX1 : OUT STD_LOGIC;
        HEX2 : OUT STD_LOGIC;
        HEX3 : OUT STD_LOGIC;
        HEX4 : OUT STD_LOGIC;
        HEX5 : OUT STD_LOGIC;
        HEX6 : OUT STD_LOGIC;
        HEX7 : OUT STD_LOGIC;
        HEX21 : OUT STD_LOGIC;
        HEX22 : OUT STD_LOGIC;
        HEX23 : OUT STD_LOGIC;
        HEX24 : OUT STD_LOGIC;
        HEX25 : OUT STD_LOGIC;
        HEX26 : OUT STD_LOGIC;
        HEX27 : OUT STD_LOGIC;
        Validation : OUT STD_LOGIC
    );
END AffichagePorte;

ARCHITECTURE BEHAVIOR OF AffichagePorte IS
    TYPE type_fstate IS (ferme,SEMIOUVERT,OUVERT);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,X)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ferme;
            HEX1 <= '0';
            HEX2 <= '0';
            HEX3 <= '0';
            HEX4 <= '0';
            HEX5 <= '0';
            HEX6 <= '0';
            HEX7 <= '0';
            HEX21 <= '0';
            HEX22 <= '0';
            HEX23 <= '0';
            HEX24 <= '0';
            HEX25 <= '0';
            HEX26 <= '0';
            HEX27 <= '0';
            Validation <= '0';
        ELSE
            HEX1 <= '0';
            HEX2 <= '0';
            HEX3 <= '0';
            HEX4 <= '0';
            HEX5 <= '0';
            HEX6 <= '0';
            HEX7 <= '0';
            HEX21 <= '0';
            HEX22 <= '0';
            HEX23 <= '0';
            HEX24 <= '0';
            HEX25 <= '0';
            HEX26 <= '0';
            HEX27 <= '0';
            Validation <= '0';
            CASE fstate IS
                WHEN ferme =>
                    IF (NOT((X = '1'))) THEN
                        reg_fstate <= SEMIOUVERT;
                    ELSIF ((X = '1')) THEN
                        reg_fstate <= ferme;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ferme;
                    END IF;

                    HEX5 <= '0';

                    HEX4 <= '0';

                    HEX6 <= '0';

                    HEX24 <= '0';

                    HEX1 <= '0';

                    HEX2 <= '0';

                    HEX25 <= '0';

                    HEX7 <= '1';

                    HEX3 <= '0';

                    Validation <= '1';

                    HEX26 <= '0';

                    HEX21 <= '0';

                    HEX27 <= '1';

                    HEX23 <= '0';

                    HEX22 <= '0';
                WHEN SEMIOUVERT =>
                    IF ((X = '1')) THEN
                        reg_fstate <= ferme;
                    ELSIF (NOT((X = '1'))) THEN
                        reg_fstate <= OUVERT;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SEMIOUVERT;
                    END IF;

                    HEX5 <= '1';

                    HEX4 <= '0';

                    HEX6 <= '1';

                    HEX24 <= '0';

                    HEX1 <= '0';

                    HEX2 <= '0';

                    HEX25 <= '0';

                    HEX7 <= '1';

                    HEX3 <= '0';

                    Validation <= '0';

                    HEX26 <= '0';

                    HEX21 <= '0';

                    HEX27 <= '1';

                    HEX23 <= '1';

                    HEX22 <= '1';
                WHEN OUVERT =>
                    IF ((X = '1')) THEN
                        reg_fstate <= SEMIOUVERT;
                    ELSIF (NOT((X = '1'))) THEN
                        reg_fstate <= OUVERT;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= OUVERT;
                    END IF;

                    HEX5 <= '1';

                    HEX4 <= '1';

                    HEX6 <= '1';

                    HEX24 <= '1';

                    HEX1 <= '1';

                    HEX2 <= '0';

                    HEX25 <= '0';

                    HEX7 <= '1';

                    HEX3 <= '0';

                    Validation <= '0';

                    HEX26 <= '0';

                    HEX21 <= '1';

                    HEX27 <= '1';

                    HEX23 <= '1';

                    HEX22 <= '1';
                WHEN OTHERS => 
                    HEX1 <= 'X';
                    HEX2 <= 'X';
                    HEX3 <= 'X';
                    HEX4 <= 'X';
                    HEX5 <= 'X';
                    HEX6 <= 'X';
                    HEX7 <= 'X';
                    HEX21 <= 'X';
                    HEX22 <= 'X';
                    HEX23 <= 'X';
                    HEX24 <= 'X';
                    HEX25 <= 'X';
                    HEX26 <= 'X';
                    HEX27 <= 'X';
                    Validation <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
