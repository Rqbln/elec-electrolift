-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Thu Nov  2 17:50:43 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY AlarMaintenance IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Maintenance : IN STD_LOGIC := '0';
        Alarme : IN STD_LOGIC := '0';
        buzzer : OUT STD_LOGIC;
        outAlarme : OUT STD_LOGIC;
        freezeAscenseur : OUT STD_LOGIC;
        outMaintenance : OUT STD_LOGIC
    );
END AlarMaintenance;

ARCHITECTURE BEHAVIOR OF AlarMaintenance IS
    TYPE type_fstate IS (state1,state2,state3,state4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Maintenance,Alarme)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            buzzer <= '0';
            outAlarme <= '0';
            freezeAscenseur <= '0';
            outMaintenance <= '0';
        ELSE
            buzzer <= '0';
            outAlarme <= '0';
            freezeAscenseur <= '0';
            outMaintenance <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((NOT((Maintenance = '1')) AND (Alarme = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF (((Maintenance = '1') AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state2;
                    ELSIF (((Maintenance = '1') AND (Alarme = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF ((NOT((Maintenance = '1')) AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    buzzer <= '0';

                    outMaintenance <= '0';

                    outAlarme <= '0';

                    freezeAscenseur <= '0';
                WHEN state2 =>
                    IF ((NOT((Maintenance = '1')) AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((Maintenance = '1') AND (Alarme = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF ((NOT((Maintenance = '1')) AND (Alarme = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF (((Maintenance = '1') AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    buzzer <= '0';

                    outMaintenance <= '1';

                    outAlarme <= '0';

                    freezeAscenseur <= '1';
                WHEN state3 =>
                    IF ((NOT((Maintenance = '1')) AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((Maintenance = '1') AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state2;
                    ELSIF (((Maintenance = '1') AND (Alarme = '1'))) THEN
                        reg_fstate <= state4;
                    ELSIF ((NOT((Maintenance = '1')) AND (Alarme = '1'))) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    buzzer <= '1';

                    outMaintenance <= '0';

                    outAlarme <= '1';

                    freezeAscenseur <= '1';
                WHEN state4 =>
                    IF ((NOT((Maintenance = '1')) AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((Maintenance = '1') AND NOT((Alarme = '1')))) THEN
                        reg_fstate <= state2;
                    ELSIF ((NOT((Maintenance = '1')) AND (Alarme = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF (((Maintenance = '1') AND (Alarme = '1'))) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    buzzer <= '0';

                    outMaintenance <= '0';

                    outAlarme <= '0';

                    freezeAscenseur <= '0';
                WHEN OTHERS => 
                    buzzer <= 'X';
                    outAlarme <= 'X';
                    freezeAscenseur <= 'X';
                    outMaintenance <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
