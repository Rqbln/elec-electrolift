-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Fri Oct 27 14:14:54 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PRESIDENT IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        KEY0 : IN STD_LOGIC := '0';
        KEY1 : IN STD_LOGIC := '0';
        Z : OUT STD_LOGIC
    );
END PRESIDENT;

ARCHITECTURE BEHAVIOR OF PRESIDENT IS
    TYPE type_fstate IS (state2,state4,state5,state6,state7,state3,state1,state8,state9,state10,state11,state12);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,KEY0,KEY1)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            Z <= '0';
        ELSE
            Z <= '0';
            CASE fstate IS
                WHEN state2 =>
                    IF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state2;
                    ELSIF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;
                WHEN state4 =>
                    IF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state4;
                    ELSIF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;
                WHEN state5 =>
                    IF ((NOT((KEY1 = '1')) AND NOT((KEY0 = '1')))) THEN
                        reg_fstate <= state5;
                    ELSIF (((KEY1 = '1') AND NOT((KEY0 = '1')))) THEN
                        reg_fstate <= state6;
                    ELSIF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;
                WHEN state6 =>
                    IF (((KEY1 = '1') AND NOT((KEY0 = '1')))) THEN
                        reg_fstate <= state6;
                    ELSIF ((NOT((KEY1 = '1')) AND NOT((KEY0 = '1')))) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;
                WHEN state7 =>
                    IF ((NOT((KEY1 = '1')) AND NOT((KEY0 = '1')))) THEN
                        reg_fstate <= state7;
                    ELSIF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state8;
                    ELSIF ((NOT((KEY0 = '1')) AND (KEY1 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;
                WHEN state3 =>
                    IF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state3;
                    ELSIF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state4;
                    ELSIF ((NOT((KEY0 = '1')) AND (KEY1 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;
                WHEN state1 =>
                    IF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;
                WHEN state8 =>
                    IF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state8;
                    ELSIF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;
                WHEN state9 =>
                    IF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state9;
                    ELSIF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state10;
                    ELSIF ((NOT((KEY0 = '1')) AND (KEY1 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;
                WHEN state10 =>
                    IF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state10;
                    ELSIF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state11;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;
                WHEN state11 =>
                    IF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state12;
                    ELSIF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state11;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state11;
                    END IF;

                    Z <= '1';
                WHEN state12 =>
                    IF ((NOT((KEY0 = '1')) AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((KEY0 = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state12;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state12;
                    END IF;

                    Z <= '0';
                WHEN OTHERS => 
                    Z <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
