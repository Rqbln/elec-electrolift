-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
-- CREATED		"Tue Oct 10 16:54:20 2023"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY DivHorlogemodif IS 
	PORT
	(
		CLOCK_50Mhz :  IN  STD_LOGIC;
		LEDR0 :  OUT  STD_LOGIC;
		LEDR1 :  OUT  STD_LOGIC;
		LEDR2 :  OUT  STD_LOGIC;
		LEDR3 :  OUT  STD_LOGIC;
		LEDR4 :  OUT  STD_LOGIC;
		LEDR5 :  OUT  STD_LOGIC;
		LEDR6 :  OUT  STD_LOGIC;
		LEDR7 :  OUT  STD_LOGIC;
		LEDR8 :  OUT  STD_LOGIC;
		LEDR9 :  OUT  STD_LOGIC
	);
END DivHorlogemodif;

ARCHITECTURE bdf_type OF DivHorlogemodif IS 

COMPONENT my_74390a
	PORT(CLKB1 : IN STD_LOGIC;
		 CLKA1 : IN STD_LOGIC;
		 CLR1 : IN STD_LOGIC;
		 CLKB2 : IN STD_LOGIC;
		 CLKA2 : IN STD_LOGIC;
		 CLR2 : IN STD_LOGIC;
		 QD11 : OUT STD_LOGIC;
		 QC11 : OUT STD_LOGIC;
		 QB11 : OUT STD_LOGIC;
		 QA11 : OUT STD_LOGIC;
		 QD22 : OUT STD_LOGIC;
		 QC22 : OUT STD_LOGIC;
		 QB22 : OUT STD_LOGIC;
		 QA22 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT my_7490
	PORT(SET9A : IN STD_LOGIC;
		 SET9B : IN STD_LOGIC;
		 CLRA : IN STD_LOGIC;
		 CLRB : IN STD_LOGIC;
		 CLKA : IN STD_LOGIC;
		 CLKB : IN STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC;
		 QD : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;


BEGIN 
LEDR9 <= CLOCK_50Mhz;
LEDR0 <= SYNTHESIZED_WIRE_40;
LEDR1 <= SYNTHESIZED_WIRE_40;
LEDR2 <= SYNTHESIZED_WIRE_40;
LEDR3 <= SYNTHESIZED_WIRE_40;
LEDR4 <= SYNTHESIZED_WIRE_40;
LEDR5 <= SYNTHESIZED_WIRE_40;
LEDR6 <= SYNTHESIZED_WIRE_40;
SYNTHESIZED_WIRE_35 <= '0';
SYNTHESIZED_WIRE_36 <= '0';
SYNTHESIZED_WIRE_37 <= '0';
SYNTHESIZED_WIRE_38 <= '0';
SYNTHESIZED_WIRE_39 <= '0';



b2v_inst1 : my_74390a
PORT MAP(CLKB1 => CLOCK_50Mhz,
		 CLKA1 => SYNTHESIZED_WIRE_0,
		 CLR1 => SYNTHESIZED_WIRE_35,
		 CLKB2 => SYNTHESIZED_WIRE_2,
		 CLKA2 => SYNTHESIZED_WIRE_3,
		 CLR2 => SYNTHESIZED_WIRE_35,
		 QD11 => SYNTHESIZED_WIRE_0,
		 QA11 => SYNTHESIZED_WIRE_2,
		 QD22 => SYNTHESIZED_WIRE_3,
		 QA22 => SYNTHESIZED_WIRE_11);





b2v_inst14 : my_74390a
PORT MAP(CLKB1 => SYNTHESIZED_WIRE_5,
		 CLKA1 => SYNTHESIZED_WIRE_6,
		 CLR1 => SYNTHESIZED_WIRE_36,
		 CLKB2 => SYNTHESIZED_WIRE_8,
		 CLKA2 => SYNTHESIZED_WIRE_9,
		 CLR2 => SYNTHESIZED_WIRE_36,
		 QD11 => SYNTHESIZED_WIRE_6,
		 QA11 => SYNTHESIZED_WIRE_8,
		 QD22 => SYNTHESIZED_WIRE_9,
		 QA22 => SYNTHESIZED_WIRE_22);




b2v_inst7 : my_74390a
PORT MAP(CLKB1 => SYNTHESIZED_WIRE_11,
		 CLKA1 => SYNTHESIZED_WIRE_12,
		 CLR1 => SYNTHESIZED_WIRE_37,
		 CLKB2 => SYNTHESIZED_WIRE_14,
		 CLKA2 => SYNTHESIZED_WIRE_15,
		 CLR2 => SYNTHESIZED_WIRE_37,
		 QD11 => SYNTHESIZED_WIRE_12,
		 QA11 => SYNTHESIZED_WIRE_14,
		 QD22 => SYNTHESIZED_WIRE_15,
		 QA22 => SYNTHESIZED_WIRE_5);


b2v_inst8 : my_7490
PORT MAP(SET9A => SYNTHESIZED_WIRE_38,
		 SET9B => SYNTHESIZED_WIRE_38,
		 CLRA => SYNTHESIZED_WIRE_38,
		 CLRB => SYNTHESIZED_WIRE_38,
		 CLKA => SYNTHESIZED_WIRE_21,
		 CLKB => SYNTHESIZED_WIRE_22,
		 QA => SYNTHESIZED_WIRE_28,
		 QD => SYNTHESIZED_WIRE_21);


b2v_inst9 : my_7490
PORT MAP(SET9A => SYNTHESIZED_WIRE_39,
		 SET9B => SYNTHESIZED_WIRE_39,
		 CLRA => SYNTHESIZED_WIRE_39,
		 CLRB => SYNTHESIZED_WIRE_39,
		 CLKA => SYNTHESIZED_WIRE_39,
		 CLKB => SYNTHESIZED_WIRE_28,
		 QA => LEDR8,
		 QB => LEDR7,
		 QD => SYNTHESIZED_WIRE_40);


END bdf_type;