-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Sat Nov  4 14:54:16 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY AlarmeClock IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        divHorloge : IN STD_LOGIC := '0';
        KEY1 : IN STD_LOGIC := '0';
        output1 : OUT STD_LOGIC
    );
END AlarmeClock;

ARCHITECTURE BEHAVIOR OF AlarmeClock IS
    TYPE type_fstate IS (state1,state2,state3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,divHorloge,KEY1)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            output1 <= '0';
        ELSE
            output1 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF (((divHorloge = '1') AND (KEY1 = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF ((NOT((divHorloge = '1')) AND (KEY1 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    output1 <= '0';
                WHEN state2 =>
                    IF (((divHorloge = '1') AND NOT((KEY1 = '1')))) THEN
                        reg_fstate <= state2;
                    ELSIF ((KEY1 = '1')) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    output1 <= '1';
                WHEN state3 =>
                    IF (NOT((KEY1 = '1'))) THEN
                        reg_fstate <= state2;
                    ELSIF ((KEY1 = '1')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    output1 <= '1';
                WHEN OTHERS => 
                    output1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
