-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Sat Oct 28 11:11:48 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY moving_zebitest2 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        sw0 : IN STD_LOGIC := '0';
        sw1 : IN STD_LOGIC := '0';
        sw2 : IN STD_LOGIC := '0';
        led0 : OUT STD_LOGIC;
        led1 : OUT STD_LOGIC;
        led2 : OUT STD_LOGIC
    );
END moving_zebitest2;

ARCHITECTURE BEHAVIOR OF moving_zebitest2 IS
    TYPE type_fstate IS (RDC,E1,E2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sw0,sw1,sw2)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= RDC;
            led0 <= '0';
            led1 <= '0';
            led2 <= '0';
        ELSE
            led0 <= '0';
            led1 <= '0';
            led2 <= '0';
            CASE fstate IS
                WHEN RDC =>
                    IF ((NOT((sw0 = '1')) AND ((sw1 = '1') OR (sw2 = '1')))) THEN
                        reg_fstate <= E1;
                    ELSIF ((sw0 = '1')) THEN
                        reg_fstate <= RDC;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= RDC;
                    END IF;

                    led2 <= '0';

                    led1 <= '0';

                    led0 <= '1';
                WHEN E1 =>
                    IF (((sw0 = '1') AND (NOT((sw1 = '1')) AND NOT((sw2 = '1'))))) THEN
                        reg_fstate <= RDC;
                    ELSIF ((NOT((sw1 = '1')) AND (sw2 = '1'))) THEN
                        reg_fstate <= E2;
                    ELSIF ((sw1 = '1')) THEN
                        reg_fstate <= E1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E1;
                    END IF;

                    led2 <= '0';

                    led1 <= '1';

                    led0 <= '0';
                WHEN E2 =>
                    IF ((NOT((sw2 = '1')) AND ((sw1 = '1') OR (sw0 = '1')))) THEN
                        reg_fstate <= E1;
                    ELSIF ((sw2 = '1')) THEN
                        reg_fstate <= E2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E2;
                    END IF;

                    led2 <= '1';

                    led1 <= '0';

                    led0 <= '0';
                WHEN OTHERS => 
                    led0 <= 'X';
                    led1 <= 'X';
                    led2 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
