-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
-- CREATED		"Tue Oct 10 15:07:48 2023"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY my_74390A IS 
	PORT
	(
		CLKB1 :  IN  STD_LOGIC;
		CLKA1 :  IN  STD_LOGIC;
		CLR1 :  IN  STD_LOGIC;
		CLKB2 :  IN  STD_LOGIC;
		CLKA2 :  IN  STD_LOGIC;
		CLR2 :  IN  STD_LOGIC;
		QD11 :  OUT  STD_LOGIC;
		QC11 :  OUT  STD_LOGIC;
		QB11 :  OUT  STD_LOGIC;
		QA11 :  OUT  STD_LOGIC;
		QD22 :  OUT  STD_LOGIC;
		QC22 :  OUT  STD_LOGIC;
		QB22 :  OUT  STD_LOGIC;
		QA22 :  OUT  STD_LOGIC
	);
END my_74390A;

ARCHITECTURE bdf_type OF my_74390A IS 

SIGNAL	QA11_INTERNAL :  STD_LOGIC;
SIGNAL	QB11_INTERNAL :  STD_LOGIC;
SIGNAL	QC11_INTERNAL :  STD_LOGIC;
SIGNAL	QD11_INTERNAL :  STD_LOGIC;
SIGNAL	QA22_INTERNAL :  STD_LOGIC;
SIGNAL	QB22_INTERNAL :  STD_LOGIC;
SIGNAL	QC22_INTERNAL :  STD_LOGIC;
SIGNAL	QD22_INTERNAL :  STD_LOGIC;
SIGNAL	QB_ALTERA_SYNTHESIZED1 :  STD_LOGIC;
SIGNAL	QB_ALTERA_SYNTHESIZED2 :  STD_LOGIC;
SIGNAL	QC_ALTERA_SYNTHESIZED1 :  STD_LOGIC;
SIGNAL	QC_ALTERA_SYNTHESIZED2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_35 <= '1';




SYNTHESIZED_WIRE_25 <= NOT(QB11_INTERNAL);



SYNTHESIZED_WIRE_5 <= NOT(CLKB1);



SYNTHESIZED_WIRE_29 <= NOT(SYNTHESIZED_WIRE_0 AND CLKB1);


SYNTHESIZED_WIRE_0 <= NOT(QD11_INTERNAL);



SYNTHESIZED_WIRE_34 <= NOT(CLR1);



SYNTHESIZED_WIRE_33 <= NOT(CLKA1);



SYNTHESIZED_WIRE_21 <= NOT(CLKA2);



SYNTHESIZED_WIRE_36 <= NOT(CLR2);



SYNTHESIZED_WIRE_1 <= NOT(QD22_INTERNAL);



SYNTHESIZED_WIRE_9 <= NOT(CLKB2);



SYNTHESIZED_WIRE_13 <= NOT(QB22_INTERNAL);



SYNTHESIZED_WIRE_17 <= NOT(SYNTHESIZED_WIRE_1 AND CLKB2);


PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_34)
VARIABLE synthesized_var_for_1QD : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	synthesized_var_for_1QD := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_5)) THEN
	synthesized_var_for_1QD := (NOT(synthesized_var_for_1QD) AND SYNTHESIZED_WIRE_4) OR (synthesized_var_for_1QD AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QD11_INTERNAL <= synthesized_var_for_1QD;
END PROCESS;


SYNTHESIZED_WIRE_8 <= QC_ALTERA_SYNTHESIZED2 AND QB_ALTERA_SYNTHESIZED2;


PROCESS(SYNTHESIZED_WIRE_9,SYNTHESIZED_WIRE_36)
VARIABLE synthesized_var_for_2QD : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_36 = '0') THEN
	synthesized_var_for_2QD := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_9)) THEN
	synthesized_var_for_2QD := (NOT(synthesized_var_for_2QD) AND SYNTHESIZED_WIRE_8) OR (synthesized_var_for_2QD AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QD22_INTERNAL <= synthesized_var_for_2QD;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_13,SYNTHESIZED_WIRE_36)
VARIABLE synthesized_var_for_2QC : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_36 = '0') THEN
	synthesized_var_for_2QC := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_13)) THEN
	synthesized_var_for_2QC := (NOT(synthesized_var_for_2QC) AND SYNTHESIZED_WIRE_35) OR (synthesized_var_for_2QC AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QC22_INTERNAL <= synthesized_var_for_2QC;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_17,SYNTHESIZED_WIRE_36)
VARIABLE synthesized_var_for_2QB : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_36 = '0') THEN
	synthesized_var_for_2QB := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_17)) THEN
	synthesized_var_for_2QB := (NOT(synthesized_var_for_2QB) AND SYNTHESIZED_WIRE_35) OR (synthesized_var_for_2QB AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QB22_INTERNAL <= synthesized_var_for_2QB;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_21,SYNTHESIZED_WIRE_36)
VARIABLE synthesized_var_for_2QA : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_36 = '0') THEN
	synthesized_var_for_2QA := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_21)) THEN
	synthesized_var_for_2QA := (NOT(synthesized_var_for_2QA) AND SYNTHESIZED_WIRE_35) OR (synthesized_var_for_2QA AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QA22_INTERNAL <= synthesized_var_for_2QA;
END PROCESS;


SYNTHESIZED_WIRE_4 <= QC_ALTERA_SYNTHESIZED1 AND QB_ALTERA_SYNTHESIZED1;


PROCESS(SYNTHESIZED_WIRE_25,SYNTHESIZED_WIRE_34)
VARIABLE synthesized_var_for_1QC : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	synthesized_var_for_1QC := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_25)) THEN
	synthesized_var_for_1QC := (NOT(synthesized_var_for_1QC) AND SYNTHESIZED_WIRE_35) OR (synthesized_var_for_1QC AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QC11_INTERNAL <= synthesized_var_for_1QC;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_29,SYNTHESIZED_WIRE_34)
VARIABLE synthesized_var_for_1QB : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	synthesized_var_for_1QB := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_29)) THEN
	synthesized_var_for_1QB := (NOT(synthesized_var_for_1QB) AND SYNTHESIZED_WIRE_35) OR (synthesized_var_for_1QB AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QB11_INTERNAL <= synthesized_var_for_1QB;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_33,SYNTHESIZED_WIRE_34)
VARIABLE synthesized_var_for_1QA : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_34 = '0') THEN
	synthesized_var_for_1QA := '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_33)) THEN
	synthesized_var_for_1QA := (NOT(synthesized_var_for_1QA) AND SYNTHESIZED_WIRE_35) OR (synthesized_var_for_1QA AND (NOT(SYNTHESIZED_WIRE_35)));
END IF;
	QA11_INTERNAL <= synthesized_var_for_1QA;
END PROCESS;

QC_ALTERA_SYNTHESIZED1 <= QC11_INTERNAL;
QB_ALTERA_SYNTHESIZED1 <= QB11_INTERNAL;
QC_ALTERA_SYNTHESIZED2 <= QC22_INTERNAL;
QB_ALTERA_SYNTHESIZED2 <= QB22_INTERNAL;
QD11 <= QD11_INTERNAL;
QC11 <= QC_ALTERA_SYNTHESIZED1;
QB11 <= QB_ALTERA_SYNTHESIZED1;
QA11 <= QA11_INTERNAL;
QD22 <= QD22_INTERNAL;
QC22 <= QC_ALTERA_SYNTHESIZED2;
QB22 <= QB_ALTERA_SYNTHESIZED2;
QA22 <= QA22_INTERNAL;

END bdf_type;